module design_example(
  output bit [7:0] addr
);
  initial addr <= 10;
endmodule
