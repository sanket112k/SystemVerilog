//environment
