program design_example(
  output reg [7:0] addr
);
  initial addr <= 10;
endprogram
