interface intf();
  logic a;
  logic b;
  logic c;
  logic sum;
  logic cout;
  
  //clocking block
  //modport
endinterface
