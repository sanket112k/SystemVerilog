program testbench(
  input reg [7:0] addr
);
  initial $display("\t Addr = %0d", addr);
endprogram
