//scoreboard
