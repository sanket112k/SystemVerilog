interface intf(
  input bit clk
);
  logic reset;
  logic data;
  logic q;
  
  // clocking block
  // modport
  
endinterface
